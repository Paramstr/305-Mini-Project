LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY ball IS
    PORT
        ( clk                       : IN std_logic;
          pixel_row, pixel_column    : IN std_logic_vector(9 DOWNTO 0);
          red, green, blue           : OUT std_logic);       
END ball;

architecture behavior of ball is

SIGNAL ball_on                   : std_logic;
SIGNAL size                      : std_logic_vector(9 DOWNTO 0);  
SIGNAL ball_x_pos,ball_y_pos    : std_logic_vector(9 DOWNTO 0);





BEGIN           

size <= CONV_STD_LOGIC_VECTOR(8,10); -- Size of the main body
-- ball_x_pos and ball_y_pos show the (x,y) for the centre of ball
ball_x_pos <= CONV_STD_LOGIC_VECTOR(128,10);
ball_y_pos <= CONV_STD_LOGIC_VECTOR(240,10);



ball_on <= '1' when ( ('0' & ball_x_pos <= '0' & pixel_column + size) and ('0' & pixel_column <= '0' & ball_x_pos + size) 	-- x_pos - size <= pixel_column <= x_pos + size
 					and ('0' & ball_y_pos <= pixel_row + size) and ('0' & pixel_row <= ball_y_pos + size) )  else	-- y_pos - size <= pixel_row <= y_pos + size
 			'0';



-- Colours for pixel data on video signal
-- Keeping background white and square in red
Red <=  '1';
-- Turn off Green and Blue when displaying square
Green <= not ball_on;
Blue <=  not ball_on;

END behavior;

